module main

// $ v -b wasm hello_world.v
// $ wasmer hello_world.wasm
// Hello WASI!
//

fn main() {
	println('Hello WASI!')
	println('Hello WASI!')
}
